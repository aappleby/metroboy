`include "types.sv"

import types::*;

module CPU(input bool x);
endmodule;