//--------------------------------------------------------------------------------
// MODULE:       uart_hello
// MODULEPARAMS: 
// INPUTS:       i_cts, i_idle, 
// OUTPUTS:      o_data, o_req, o_done, 
// LOCALPARAMS:  message_len, cursor_bits, 
// FIELDS:       state, cursor, memory, data, 
// SUBMODULES:   
// TASKS:        
// FUNCTIONS:    
/* verilator lint_off WIDTH */
`default_nettype none

`include "metron.h.sv"

//==============================================================================

module uart_hello
(clk, rst_n, i_cts, i_idle, o_data, o_req, o_done);
  /*verilator public_module*/
  
  input logic clk;
  input logic rst_n;
  input bool i_cts;
  input bool i_idle; 

  localparam int message_len = 'd512;
  localparam int cursor_bits = $clog2(message_len);

  typedef enum { WAIT, SEND, DONE } e_state;
  logic[1:0] state;
  logic[cursor_bits-1:0] cursor;
  logic[7:0] memory['d512];
  logic[7:0] data;

  output logic[7:0] o_data;
  output logic o_req;
  output logic o_done;

  //----------------------------------------

  initial begin : INIT
    $readmemh("obj/message.hex", memory, 'd0, 'd511);
    o_data = 'd0;
    o_req = 'd0;
    o_done = 'd0;
  end

  //----------------------------------------

  always_ff @(posedge clk, negedge rst_n) begin : TICK
    if (!rst_n) begin
      state <= WAIT;
      cursor <= 'd0;
    end
    else begin
      data <= memory[cursor];
      if (state == WAIT && i_idle) begin
        state <= SEND;
      end
      else if (state == SEND && i_cts) begin
        if (cursor == (message_len - 'd1)) state <= DONE;
        cursor <= cursor + 'd1;
      end
      else if (state == DONE) begin
        //state = WAIT;
        cursor <= 'd0;
      end
    end
  end

  //----------------------------------------

  always_comb begin : TOCK
    o_data = data;
    o_req = state == SEND;
    o_done = state == DONE;
  end

endmodule

//==============================================================================
